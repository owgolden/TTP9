`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

  // // Data inputs
  //  wire [11:0] in;
  //  assign ui_in[0]  = in[0];
  //  assign ui_in[1]  = in[1];
  //  assign ui_in[2]  = in[2];
  //  assign ui_in[3]  = in[3];
  //  assign ui_in[4]  = in[4];
  //  assign ui_in[5]  = in[5];
  //  assign ui_in[6]  = in[6];
  //  assign ui_in[7]  = in[7];
  //  assign uio_in[0] = in[8];
  //  assign uio_in[1] = in[9];
  //  assign uio_in[2] = in[10];
  //  assign uio_in[3] = in[11];

  //  // input for selecting the register ( "0" - duty_reg, "1" - period_reg)
  //  wire sel;
  //  assign uio_in[6] = sel;

  //  // input for write enable ("0" - do nothing,"1" - write selected register)
  //  wire wr_en;
  //  assign uio_in[7] = wr_en;

  //  // PWM output 
  //  wire pwm_out;
  //  assign uo_out[0] = pwm_out;
   
  // Replace tt_um_example with your module name:
  tt_um_samuelm_pwm_generator user_project(

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(1'b1),
      .VGND(1'b0),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
